module mimas (gpio);

output [31:0] gpio;

wire [31:0] gpio;

assign gpio = 8'hAAAAAAAA;

endmodule
